netcdf lis_input {
dimensions:
	east_west = 1440 ;
	north_south = 600 ;
	east_west_b = 1444 ;
	north_south_b = 604 ;
	east_west_GDAS_T126 = 384 ;
	north_south_GDAS_T126 = 190 ;
	east_west_GDAS_T170 = 512 ;
	north_south_GDAS_T170 = 256 ;
	east_west_GDAS_T254 = 768 ;
	north_south_GDAS_T254 = 384 ;
	east_west_GDAS_T382 = 1152 ;
	north_south_GDAS_T382 = 576 ;
	east_west_GDAS_T574 = 1760 ;
	north_south_GDAS_T574 = 880 ;
	east_west_GDAS_T1534 = 3072 ;
	north_south_GDAS_T1534 = 1536 ;
	month = 12 ;
	time = 1 ;
	sfctypes = 20 ;
	soiltypes = 16 ;
	elevbins = 1 ;
variables:
	float time(time) ;
	float LANDMASK(north_south, east_west) ;
		LANDMASK:standard_name = "LANDMASK" ;
		LANDMASK:units = "" ;
		LANDMASK:scale_factor = 1.f ;
		LANDMASK:add_offset = 0.f ;
		LANDMASK:missing_value = -9999.f ;
		LANDMASK:vmin = 0.f ;
		LANDMASK:vmax = 0.f ;
		LANDMASK:num_bins = 1 ;
	float SURFACETYPE(sfctypes, north_south, east_west) ;
		SURFACETYPE:standard_name = "Surface type" ;
		SURFACETYPE:units = "-" ;
		SURFACETYPE:scale_factor = 1.f ;
		SURFACETYPE:add_offset = 0.f ;
		SURFACETYPE:missing_value = -9999.f ;
		SURFACETYPE:vmin = 0.f ;
		SURFACETYPE:vmax = 0.f ;
		SURFACETYPE:num_bins = 20 ;
	float LANDCOVER(sfctypes, north_south, east_west) ;
		LANDCOVER:standard_name = "MODIS-IGBP (NCEP-modified) landcover map" ;
		LANDCOVER:units = "" ;
		LANDCOVER:scale_factor = 1.f ;
		LANDCOVER:add_offset = 0.f ;
		LANDCOVER:missing_value = -9999.f ;
		LANDCOVER:vmin = 0.f ;
		LANDCOVER:vmax = 0.f ;
		LANDCOVER:num_bins = 20 ;
	float TEXTURE(soiltypes, north_south, east_west) ;
		TEXTURE:standard_name = "(NCAR) STATSGO+FAO blended soil texture map" ;
		TEXTURE:units = "" ;
		TEXTURE:scale_factor = 1.f ;
		TEXTURE:add_offset = 0.f ;
		TEXTURE:missing_value = -9999.f ;
		TEXTURE:vmin = 0.f ;
		TEXTURE:vmax = 0.f ;
		TEXTURE:num_bins = 16 ;
	float ELEVFGRD(north_south, east_west) ;
		ELEVFGRD:standard_name = "Elevation Area Fraction" ;
		ELEVFGRD:units = "-" ;
		ELEVFGRD:scale_factor = 1.f ;
		ELEVFGRD:add_offset = 0.f ;
		ELEVFGRD:missing_value = -9999.f ;
		ELEVFGRD:vmin = 0.f ;
		ELEVFGRD:vmax = 0.f ;
		ELEVFGRD:num_bins = 1 ;
	float ELEVATION(north_south, east_west) ;
		ELEVATION:standard_name = "SRTM (Native) elevation" ;
		ELEVATION:units = "m" ;
		ELEVATION:scale_factor = 1.f ;
		ELEVATION:add_offset = 0.f ;
		ELEVATION:missing_value = -9999.f ;
		ELEVATION:vmin = 0.f ;
		ELEVATION:vmax = 0.f ;
		ELEVATION:num_bins = 1 ;
	float GREENNESS(month, north_south, east_west) ;
		GREENNESS:standard_name = "NCEP (Native) monthly greenness fraction climatology" ;
		GREENNESS:units = "-" ;
		GREENNESS:scale_factor = 1.f ;
		GREENNESS:add_offset = 0.f ;
		GREENNESS:missing_value = -9999.f ;
		GREENNESS:vmin = 0.f ;
		GREENNESS:vmax = 0.f ;
		GREENNESS:num_bins = 1 ;
	float SHDMIN(north_south, east_west) ;
		SHDMIN:standard_name = "NCEP (Native) min greenness" ;
		SHDMIN:units = "-" ;
		SHDMIN:scale_factor = 1.f ;
		SHDMIN:add_offset = 0.f ;
		SHDMIN:missing_value = -9999.f ;
		SHDMIN:vmin = 0.f ;
		SHDMIN:vmax = 0.f ;
		SHDMIN:num_bins = 1 ;
	float SHDMAX(north_south, east_west) ;
		SHDMAX:standard_name = "NCEP (Native) max greenness" ;
		SHDMAX:units = "-" ;
		SHDMAX:scale_factor = 1.f ;
		SHDMAX:add_offset = 0.f ;
		SHDMAX:missing_value = -9999.f ;
		SHDMAX:vmin = 0.f ;
		SHDMAX:vmax = 0.f ;
		SHDMAX:num_bins = 1 ;
	float ALBEDO(month, north_south, east_west) ;
		ALBEDO:standard_name = "NCEP (Native) monthly albedo clim" ;
		ALBEDO:units = "-" ;
		ALBEDO:scale_factor = 1.f ;
		ALBEDO:add_offset = 0.f ;
		ALBEDO:missing_value = -9999.f ;
		ALBEDO:vmin = 0.f ;
		ALBEDO:vmax = 0.f ;
		ALBEDO:num_bins = 1 ;
	float MXSNALBEDO(north_south, east_west) ;
		MXSNALBEDO:standard_name = "NCEP (Native) max snow albedo" ;
		MXSNALBEDO:units = "-" ;
		MXSNALBEDO:scale_factor = 1.f ;
		MXSNALBEDO:add_offset = 0.f ;
		MXSNALBEDO:missing_value = -9999.f ;
		MXSNALBEDO:vmin = 0.f ;
		MXSNALBEDO:vmax = 0.f ;
		MXSNALBEDO:num_bins = 1 ;
	float TBOT(north_south, east_west) ;
		TBOT:standard_name = "Noah LSM bottom temperature" ;
		TBOT:units = "K" ;
		TBOT:scale_factor = 1.f ;
		TBOT:add_offset = 0.f ;
		TBOT:missing_value = -9999.f ;
		TBOT:vmin = 0.f ;
		TBOT:vmax = 0.f ;
		TBOT:num_bins = 1 ;
	float SLOPETYPE(north_south, east_west) ;
		SLOPETYPE:standard_name = "Noah LSM slope type" ;
		SLOPETYPE:units = "-" ;
		SLOPETYPE:scale_factor = 1.f ;
		SLOPETYPE:add_offset = 0.f ;
		SLOPETYPE:missing_value = -9999.f ;
		SLOPETYPE:vmin = 0.f ;
		SLOPETYPE:vmax = 0.f ;
		SLOPETYPE:num_bins = 1 ;
	float NOAHMP36_PBLH(north_south, east_west) ;
		NOAHMP36_PBLH:standard_name = "Noah-MP LSM planetary boundary height" ;
		NOAHMP36_PBLH:units = "m" ;
		NOAHMP36_PBLH:scale_factor = 1.f ;
		NOAHMP36_PBLH:add_offset = 0.f ;
		NOAHMP36_PBLH:missing_value = -9999.f ;
		NOAHMP36_PBLH:vmin = 0.f ;
		NOAHMP36_PBLH:vmax = 0.f ;
		NOAHMP36_PBLH:num_bins = 1 ;
	float ELEV_GDAS_T126(north_south, east_west) ;
		ELEV_GDAS_T126:standard_name = "Forcing elevation for GDAS_T126" ;
		ELEV_GDAS_T126:units = "m" ;
		ELEV_GDAS_T126:scale_factor = 1.f ;
		ELEV_GDAS_T126:add_offset = 0.f ;
		ELEV_GDAS_T126:missing_value = -9999.f ;
		ELEV_GDAS_T126:vmin = 0.f ;
		ELEV_GDAS_T126:vmax = 0.f ;
		ELEV_GDAS_T126:num_bins = 1 ;
	float ELEVDIFF_GDAS_T126(north_south_GDAS_T126, east_west_GDAS_T126) ;
		ELEVDIFF_GDAS_T126:standard_name = "Forcing elevation diff for GDAS_T126" ;
		ELEVDIFF_GDAS_T126:units = "m" ;
		ELEVDIFF_GDAS_T126:scale_factor = 1.f ;
		ELEVDIFF_GDAS_T126:add_offset = 0.f ;
		ELEVDIFF_GDAS_T126:missing_value = -9999.f ;
		ELEVDIFF_GDAS_T126:vmin = 0.f ;
		ELEVDIFF_GDAS_T126:vmax = 0.f ;
		ELEVDIFF_GDAS_T126:num_bins = 1 ;
	float ELEV_GDAS_T170(north_south, east_west) ;
		ELEV_GDAS_T170:standard_name = "Forcing elevation for GDAS_T170" ;
		ELEV_GDAS_T170:units = "m" ;
		ELEV_GDAS_T170:scale_factor = 1.f ;
		ELEV_GDAS_T170:add_offset = 0.f ;
		ELEV_GDAS_T170:missing_value = -9999.f ;
		ELEV_GDAS_T170:vmin = 0.f ;
		ELEV_GDAS_T170:vmax = 0.f ;
		ELEV_GDAS_T170:num_bins = 1 ;
	float ELEVDIFF_GDAS_T170(north_south_GDAS_T170, east_west_GDAS_T170) ;
		ELEVDIFF_GDAS_T170:standard_name = "Forcing elevation diff for GDAS_T170" ;
		ELEVDIFF_GDAS_T170:units = "m" ;
		ELEVDIFF_GDAS_T170:scale_factor = 1.f ;
		ELEVDIFF_GDAS_T170:add_offset = 0.f ;
		ELEVDIFF_GDAS_T170:missing_value = -9999.f ;
		ELEVDIFF_GDAS_T170:vmin = 0.f ;
		ELEVDIFF_GDAS_T170:vmax = 0.f ;
		ELEVDIFF_GDAS_T170:num_bins = 1 ;
	float ELEV_GDAS_T254(north_south, east_west) ;
		ELEV_GDAS_T254:standard_name = "Forcing elevation for GDAS_T254" ;
		ELEV_GDAS_T254:units = "m" ;
		ELEV_GDAS_T254:scale_factor = 1.f ;
		ELEV_GDAS_T254:add_offset = 0.f ;
		ELEV_GDAS_T254:missing_value = -9999.f ;
		ELEV_GDAS_T254:vmin = 0.f ;
		ELEV_GDAS_T254:vmax = 0.f ;
		ELEV_GDAS_T254:num_bins = 1 ;
	float ELEVDIFF_GDAS_T254(north_south_GDAS_T254, east_west_GDAS_T254) ;
		ELEVDIFF_GDAS_T254:standard_name = "Forcing elevation diff for GDAS_T254" ;
		ELEVDIFF_GDAS_T254:units = "m" ;
		ELEVDIFF_GDAS_T254:scale_factor = 1.f ;
		ELEVDIFF_GDAS_T254:add_offset = 0.f ;
		ELEVDIFF_GDAS_T254:missing_value = -9999.f ;
		ELEVDIFF_GDAS_T254:vmin = 0.f ;
		ELEVDIFF_GDAS_T254:vmax = 0.f ;
		ELEVDIFF_GDAS_T254:num_bins = 1 ;
	float ELEV_GDAS_T382(north_south, east_west) ;
		ELEV_GDAS_T382:standard_name = "Forcing elevation for GDAS_T382" ;
		ELEV_GDAS_T382:units = "m" ;
		ELEV_GDAS_T382:scale_factor = 1.f ;
		ELEV_GDAS_T382:add_offset = 0.f ;
		ELEV_GDAS_T382:missing_value = -9999.f ;
		ELEV_GDAS_T382:vmin = 0.f ;
		ELEV_GDAS_T382:vmax = 0.f ;
		ELEV_GDAS_T382:num_bins = 1 ;
	float ELEVDIFF_GDAS_T382(north_south_GDAS_T382, east_west_GDAS_T382) ;
		ELEVDIFF_GDAS_T382:standard_name = "Forcing elevation diff for GDAS_T382" ;
		ELEVDIFF_GDAS_T382:units = "m" ;
		ELEVDIFF_GDAS_T382:scale_factor = 1.f ;
		ELEVDIFF_GDAS_T382:add_offset = 0.f ;
		ELEVDIFF_GDAS_T382:missing_value = -9999.f ;
		ELEVDIFF_GDAS_T382:vmin = 0.f ;
		ELEVDIFF_GDAS_T382:vmax = 0.f ;
		ELEVDIFF_GDAS_T382:num_bins = 1 ;
	float ELEV_GDAS_T574(north_south, east_west) ;
		ELEV_GDAS_T574:standard_name = "Forcing elevation for GDAS_T574" ;
		ELEV_GDAS_T574:units = "m" ;
		ELEV_GDAS_T574:scale_factor = 1.f ;
		ELEV_GDAS_T574:add_offset = 0.f ;
		ELEV_GDAS_T574:missing_value = -9999.f ;
		ELEV_GDAS_T574:vmin = 0.f ;
		ELEV_GDAS_T574:vmax = 0.f ;
		ELEV_GDAS_T574:num_bins = 1 ;
	float ELEVDIFF_GDAS_T574(north_south_GDAS_T574, east_west_GDAS_T574) ;
		ELEVDIFF_GDAS_T574:standard_name = "Forcing elevation diff for GDAS_T574" ;
		ELEVDIFF_GDAS_T574:units = "m" ;
		ELEVDIFF_GDAS_T574:scale_factor = 1.f ;
		ELEVDIFF_GDAS_T574:add_offset = 0.f ;
		ELEVDIFF_GDAS_T574:missing_value = -9999.f ;
		ELEVDIFF_GDAS_T574:vmin = 0.f ;
		ELEVDIFF_GDAS_T574:vmax = 0.f ;
		ELEVDIFF_GDAS_T574:num_bins = 1 ;
	float ELEV_GDAS_T1534(north_south, east_west) ;
		ELEV_GDAS_T1534:standard_name = "Forcing elevation for GDAS_T1534" ;
		ELEV_GDAS_T1534:units = "m" ;
		ELEV_GDAS_T1534:scale_factor = 1.f ;
		ELEV_GDAS_T1534:add_offset = 0.f ;
		ELEV_GDAS_T1534:missing_value = -9999.f ;
		ELEV_GDAS_T1534:vmin = 0.f ;
		ELEV_GDAS_T1534:vmax = 0.f ;
		ELEV_GDAS_T1534:num_bins = 1 ;
	float ELEVDIFF_GDAS_T1534(north_south_GDAS_T1534, east_west_GDAS_T1534) ;
		ELEVDIFF_GDAS_T1534:standard_name = "Forcing elevation diff for GDAS_T1534" ;
		ELEVDIFF_GDAS_T1534:units = "m" ;
		ELEVDIFF_GDAS_T1534:scale_factor = 1.f ;
		ELEVDIFF_GDAS_T1534:add_offset = 0.f ;
		ELEVDIFF_GDAS_T1534:missing_value = -9999.f ;
		ELEVDIFF_GDAS_T1534:vmin = 0.f ;
		ELEVDIFF_GDAS_T1534:vmax = 0.f ;
		ELEVDIFF_GDAS_T1534:num_bins = 1 ;
	float lat(north_south, east_west) ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.f ;
		lat:add_offset = 0.f ;
		lat:missing_value = -9999.f ;
		lat:vmin = 0.f ;
		lat:vmax = 0.f ;
	float lon(north_south, east_west) ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.f ;
		lon:add_offset = 0.f ;
		lon:missing_value = -9999.f ;
		lon:vmin = 0.f ;
		lon:vmax = 0.f ;
	float lat_b(north_south_b, east_west_b) ;
		lat_b:standard_name = "latitude_b" ;
		lat_b:units = "degrees_north" ;
		lat_b:scale_factor = 1.f ;
		lat_b:add_offset = 0.f ;
		lat_b:missing_value = -9999.f ;
		lat_b:vmin = 0.f ;
		lat_b:vmax = 0.f ;
	float lon_b(north_south_b, east_west_b) ;
		lon_b:standard_name = "longitude_b" ;
		lon_b:units = "degrees_east" ;
		lon_b:scale_factor = 1.f ;
		lon_b:add_offset = 0.f ;
		lon_b:missing_value = -9999.f ;
		lon_b:vmin = 0.f ;
		lon_b:vmax = 0.f ;

// global attributes:
		:MAP_PROJECTION = "EQUIDISTANT CYLINDRICAL" ;
		:SOUTH_WEST_CORNER_LAT = -59.875f ;
		:SOUTH_WEST_CORNER_LON = -179.875f ;
		:DX = 0.25f ;
		:DY = 0.25f ;
		:MAP_PROJECTION_GDAS_T126 = "GAUSSIAN" ;
		:NORTH_WEST_CORNER_LAT_GDAS_T126 = 89.277f ;
		:NORTH_WEST_CORNER_LON_GDAS_T126 = 0.f ;
		:SOUTH_EAST_CORNER_LAT_GDAS_T126 = -89.277f ;
		:SOUTH_EAST_CORNER_LON_GDAS_T126 = -0.938f ;
		:DI_GDAS_T126 = 0.938f ;
		:N_GDAS_T126 = 95.f ;
		:MAP_PROJECTION_GDAS_T170 = "GAUSSIAN" ;
		:NORTH_WEST_CORNER_LAT_GDAS_T170 = 89.463f ;
		:NORTH_WEST_CORNER_LON_GDAS_T170 = 0.f ;
		:SOUTH_EAST_CORNER_LAT_GDAS_T170 = -89.463f ;
		:SOUTH_EAST_CORNER_LON_GDAS_T170 = -0.703f ;
		:DI_GDAS_T170 = 0.703f ;
		:N_GDAS_T170 = 128.f ;
		:MAP_PROJECTION_GDAS_T254 = "GAUSSIAN" ;
		:NORTH_WEST_CORNER_LAT_GDAS_T254 = 89.642f ;
		:NORTH_WEST_CORNER_LON_GDAS_T254 = 0.f ;
		:SOUTH_EAST_CORNER_LAT_GDAS_T254 = -89.642f ;
		:SOUTH_EAST_CORNER_LON_GDAS_T254 = -0.469f ;
		:DI_GDAS_T254 = 0.469f ;
		:N_GDAS_T254 = 192.f ;
		:MAP_PROJECTION_GDAS_T382 = "GAUSSIAN" ;
		:NORTH_WEST_CORNER_LAT_GDAS_T382 = 89.761f ;
		:NORTH_WEST_CORNER_LON_GDAS_T382 = 0.f ;
		:SOUTH_EAST_CORNER_LAT_GDAS_T382 = -89.761f ;
		:SOUTH_EAST_CORNER_LON_GDAS_T382 = -0.313f ;
		:DI_GDAS_T382 = 0.313f ;
		:N_GDAS_T382 = 288.f ;
		:MAP_PROJECTION_GDAS_T574 = "GAUSSIAN" ;
		:NORTH_WEST_CORNER_LAT_GDAS_T574 = 89.844f ;
		:NORTH_WEST_CORNER_LON_GDAS_T574 = 0.f ;
		:SOUTH_EAST_CORNER_LAT_GDAS_T574 = -89.844f ;
		:SOUTH_EAST_CORNER_LON_GDAS_T574 = -0.205f ;
		:DI_GDAS_T574 = 0.205f ;
		:N_GDAS_T574 = 440.f ;
		:MAP_PROJECTION_GDAS_T1534 = "GAUSSIAN" ;
		:NORTH_WEST_CORNER_LAT_GDAS_T1534 = 89.91f ;
		:NORTH_WEST_CORNER_LON_GDAS_T1534 = 0.f ;
		:SOUTH_EAST_CORNER_LAT_GDAS_T1534 = -89.91f ;
		:SOUTH_EAST_CORNER_LON_GDAS_T1534 = -0.1171875f ;
		:DI_GDAS_T1534 = 0.1171875f ;
		:N_GDAS_T1534 = 768.f ;
		:INC_WATER_PTS = "false" ;
		:LANDCOVER_SCHEME = "IGBPNCEP" ;
		:NUMBER_LANDCATS = 20 ;
		:BARESOILCLASS = 16 ;
		:URBANCLASS = 13 ;
		:SNOWCLASS = 15 ;
		:WATERCLASS = 17 ;
		:WETLANDCLASS = 11 ;
		:GLACIERCLASS = 15 ;
		:NUMVEGTYPES = 17 ;
		:LANDMASK_SOURCE = "MODIS_Native" ;
		:SFCMODELS = "Noah-MP.3.6" ;
		:SOILTEXT_SCHEME = "STATSGO" ;
		:NUMBER_SOILTYPES = 19 ;
		:NUMBER_SLOPETYPES = 9 ;
		:GREENNESS_DATA_INTERVAL = "monthly" ;
		:ALBEDO_DATA_INTERVAL = "monthly" ;
		:title = "Land Data Toolkit (LDT) parameter-processed output" ;
		:institution = "NASA GSFC Hydrological Sciences Laboratory" ;
		:history = "created on date: 2015-06-19T12:01:22.281" ;
		:references = "Kumar_etal_EMS_2006, Peters-Lidard_etal_ISSE_2007" ;
		:comment = "website: http://lis.gsfc.nasa.gov/" ;
}
